module main

import vplot


